LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY half_adder IS
	PORT(
			a,b: IN STD_LOGIC;
			s, c: OUT STD_LOGIC
		);
END half_adder;
--------------------------------------------------
ARCHITECTURE behavioral OF half_adder IS
	BEGIN
		s<= a XOR b;
		c<= a AND b;
END behavioral;