LIBRARY IEEE;
USE  IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_ARITH.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;

ENTITY clk_50hz IS
		 PORT( 
		 CLK_50MHZ: IN	STD_LOGIC;
		 CLK_OUT : OUT STD_LOGIC
		 );
END clk_50hz ;
---------------------------------------------------------------

ARCHITECTURE arch OF clk_50hz IS
	SIGNAL CLK_COUNT_400HZ: STD_LOGIC_VECTOR(19 DOWNTO 0);
	SIGNAL CLK_COUNT_10HZ: STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL CLK_400HZ, CLK_10HZ : STD_LOGIC;
	BEGIN
	
	    PROCESS
			BEGIN
			 WAIT UNTIL CLK_50MHZ'EVENT AND CLK_50MHZ = '1';
						IF CLK_COUNT_400HZ < X"0F424" THEN 
						 CLK_COUNT_400HZ <= CLK_COUNT_400HZ + 1;
						ELSE
						 CLK_COUNT_400HZ <= X"00000";
						 CLK_400HZ <= NOT CLK_400HZ;
						END IF;
		END PROCESS;

		PROCESS (CLK_400HZ)
			BEGIN
				IF CLK_400HZ'EVENT AND CLK_400HZ = '1' THEN
					IF CLK_COUNT_10HZ < 19 THEN
						CLK_COUNT_10HZ <= CLK_COUNT_10HZ + 1;
					ELSE
						CLK_COUNT_10HZ <= X"00";
						CLK_10HZ <= NOT CLK_10HZ;
					END IF;
				END IF;
		END PROCESS;
		
		CLK_OUT <= CLK_10HZ;
END ARCHITECTURE;